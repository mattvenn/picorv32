`default_nettype none
/*
 *  PicoSoC - A simple example SoC using PicoRV32
 *
 *  Copyright (C) 2017  Clifford Wolf <clifford@clifford.at>
 *
 *  Permission to use, copy, modify, and/or distribute this software for any
 *  purpose with or without fee is hereby granted, provided that the above
 *  copyright notice and this permission notice appear in all copies.
 *
 *  THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 *  WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 *  MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 *  ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 *  WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 *  ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 *  OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 *
 */
module ecp5demo (
	input clk,

	output ser_tx,
	input ser_rx,
    input reset_button,

	output [7:0] leds,
    output [7:0] pmod2,

    output led1,
    output led2,

	output flash_csb,
    `ifndef SYNTH
    output flash_clk,
    `endif
	inout  flash_io0,
	inout  flash_io1,
	inout  flash_io2,
	inout  flash_io3

/*
	output debug_ser_tx,
	output debug_ser_rx,

	output debug_flash_csb,
	output debug_flash_clk,
	output debug_flash_io0,
	output debug_flash_io1,
	output debug_flash_io2,
	output debug_flash_io3
*/
);
	reg [5:0] reset_cnt = 0;
	wire resetn = &reset_cnt;

	always @(posedge clk) begin
		reset_cnt <= reset_cnt + !resetn;
        if(!reset_button) // if pressed
            reset_cnt <= 0;
	end

	wire flash_io0_oe, flash_io0_do, flash_io0_di;
	wire flash_io1_oe, flash_io1_do, flash_io1_di;
	wire flash_io2_oe, flash_io2_do, flash_io2_di;
	wire flash_io3_oe, flash_io3_do, flash_io3_di;

    `ifdef SYNTH
	wire flash_clk;
    USRMCLK u1 (.USRMCLKI(flash_clk), .USRMCLKTS(flash_csb)) /* synthesis syn_noprune=1 */;
    BBPU flash_io_buf[3:0] (
        .B({flash_io3, flash_io2, flash_io1, flash_io0}),
        .T({!flash_io3_oe,!flash_io2_oe,!flash_io1_oe, !flash_io0_oe}),
        .I({flash_io3_do, flash_io2_do, flash_io1_do, flash_io0_do}),
        .O({flash_io3_di, flash_io2_di, flash_io1_di, flash_io0_di})
    );
    `else
        // this needed for sim as ecp5 sim models not available

           SB_IO #(
                   .PIN_TYPE(6'b 1010_01),
                   .PULLUP(1'b 0)
           ) flash_io_buf [3:0] (
                   .PACKAGE_PIN({flash_io3, flash_io2, flash_io1, flash_io0}),
                   .OUTPUT_ENABLE({flash_io3_oe, flash_io2_oe, flash_io1_oe, flash_io0_oe}),
                   .D_OUT_0({flash_io3_do, flash_io2_do, flash_io1_do, flash_io0_do}),
                   .D_IN_0({flash_io3_di, flash_io2_di, flash_io1_di, flash_io0_di})
           );
    `endif

    // same address as where the gpio leds were
    wb_buttons_leds #(.BASE_ADDRESS(32'h03_00_00_00)) wb_buttons_leds_0 (
        .clk        (clk),
        .reset      (~resetn),
        .i_wb_cyc   (wbm_cyc_o),
        .i_wb_stb   (wbm_stb_o),
        .i_wb_we    (wbm_we_o),
        .i_wb_addr  (wbm_adr_o),
        .i_wb_data  (wbm_dat_o),
        .o_wb_ack   (leds_wbm_ack_i),
        .o_wb_data  (leds_wbm_dat_i),
        //.buttons    (buttons),
        .leds       (wb_leds)
    );

    user_project_wrapper  user_project_wrapper(

    // Wishbone Slave ports (WB MI A)
    .wb_clk_i       (clk),             // clock
    .wb_rst_i       (~resetn),             // reset
    .wbs_stb_i      (wbm_stb_o),            // strobe - wb_valid data
    .wbs_cyc_i      (wbm_cyc_o),            // cycle - high when during a request
    .wbs_we_i       (|wbm_we_o),             // write enable
    .wbs_sel_i      (wbm_we_o),      // which byte to read/write
    .wbs_dat_i      (wbm_dat_o),     // data in
    .wbs_adr_i      (wbm_adr_o),     // address
    .wbs_ack_o      (mph_wbm_ack_i),           // ack
    .wbs_dat_o      (mph_wbm_dat_i),    // data out

    // Logic Analyzer Signals
    .la_data_in(0),
 //   input  wire [127:0] la_data_in,
  //  output wire [127:0] la_data_out,
   // input  wire [127:0] la_oen,

    // IOs - avoid using 0-7 as they are dual purpose and maybe connected to other things
//    input  wire [`MPRJ_IO_PADS-1:0] io_in,
    .io_out(mph_io_out)
  //  output wire [`MPRJ_IO_PADS-1:0] io_oeb // active low!

    );
    wire [37:0] mph_io_out;
    assign pmod2 = mph_io_out[15:8]; // put first 8 usable outputs onto pmod2
    wire [31:0] mph_wbm_dat_i, leds_wbm_dat_i;
    wire mph_wbm_ack_i, leds_wbm_ack_i;
    assign wbm_ack_i = mph_wbm_ack_i | leds_wbm_ack_i; 
    assign wbm_dat_i = mph_wbm_dat_i | leds_wbm_dat_i; 

    wire [7:0] wb_leds;
    assign leds = wb_leds;
    assign led1 = leds[0];
    assign led2 = leds[1];
    
	localparam IDLE = 2'b00;
	localparam WBSTART = 2'b01;
	localparam WBEND = 2'b10;

	reg [1:0] state;

	wire we;
	assign we = (iomem_wstrb[0] | iomem_wstrb[1] | iomem_wstrb[2] | iomem_wstrb[3]);

	always @(posedge clk) begin
		if (~resetn) begin
			wbm_adr_o <= 0;
			wbm_dat_o <= 0;
			wbm_we_o <= 0;
			wbm_sel_o <= 0;
			wbm_stb_o <= 0;
			wbm_cyc_o <= 0;
			state <= IDLE;
		end else begin
			case (state)
				IDLE: begin
                    // wishbone is 0x0300_0000 and above
					if (iomem_valid & iomem_addr[31:24] >= 8'h03) begin
						wbm_adr_o <= iomem_addr;
						wbm_dat_o <= iomem_wdata;
						wbm_we_o <= we;
						wbm_sel_o <= iomem_wstrb;

						wbm_stb_o <= 1'b1;
						wbm_cyc_o <= 1'b1;
						state <= WBSTART;
					end else begin
						iomem_ready <= 1'b0;

						wbm_stb_o <= 1'b0;
						wbm_cyc_o <= 1'b0;
						wbm_we_o <= 1'b0;
					end
				end
				WBSTART:begin
					if (wbm_ack_i) begin
						iomem_rdata <= wbm_dat_i;
						iomem_ready <= 1'b1;

						state <= WBEND;

						wbm_stb_o <= 1'b0;
						wbm_cyc_o <= 1'b0;
						wbm_we_o <= 1'b0;
					end
				end
				WBEND: begin
					iomem_ready <= 1'b0;

					state <= IDLE;
				end
				default:
					state <= IDLE;
			endcase
		end
	end

	wire        iomem_valid;
	reg         iomem_ready;
	wire [3:0]  iomem_wstrb;
	wire [31:0] iomem_addr;
	wire [31:0] iomem_wdata;
	reg  [31:0] iomem_rdata;

    /*
	reg [31:0] gpio;
	assign leds = gpio;
    assign led1 = !gpio[0];
    assign led2 = !gpio[1];
    */

	reg [31:0] wbm_adr_o;
	reg [31:0] wbm_dat_o;
	wire [31:0] wbm_dat_i;
	reg wbm_we_o;
	reg [3:0] wbm_sel_o;
	reg wbm_stb_o;
	wire wbm_ack_i;
	reg wbm_cyc_o;

    /*
	always @(posedge clk) begin
		if (!resetn) begin
			gpio <= 0;
		end else begin
			iomem_ready <= 0;
			if (iomem_valid && !iomem_ready && iomem_addr[31:24] == 8'h 03) begin
				iomem_ready <= 1;
				iomem_rdata <= gpio;
				if (iomem_wstrb[0]) gpio[ 7: 0] <= iomem_wdata[ 7: 0];
				if (iomem_wstrb[1]) gpio[15: 8] <= iomem_wdata[15: 8];
				if (iomem_wstrb[2]) gpio[23:16] <= iomem_wdata[23:16];
				if (iomem_wstrb[3]) gpio[31:24] <= iomem_wdata[31:24];
			end
		end
	end
    */

	picosoc soc (
		.clk          (clk         ),
		.resetn       (resetn      ),
        
        .led1         (led1        ),
        .led2         (led2        ),

		.ser_tx       (ser_tx      ),
		.ser_rx       (ser_rx      ),

		.flash_csb    (flash_csb   ),
		.flash_clk    (flash_clk   ),

		.flash_io0_oe (flash_io0_oe),
		.flash_io1_oe (flash_io1_oe),
		.flash_io2_oe (flash_io2_oe),
		.flash_io3_oe (flash_io3_oe),

		.flash_io0_do (flash_io0_do),
		.flash_io1_do (flash_io1_do),
		.flash_io2_do (flash_io2_do),
		.flash_io3_do (flash_io3_do),

		.flash_io0_di (flash_io0_di),
		.flash_io1_di (flash_io1_di),
		.flash_io2_di (flash_io2_di),
		.flash_io3_di (flash_io3_di),

		.irq_5        (1'b0        ),
		.irq_6        (1'b0        ),
		.irq_7        (1'b0        ),

		.iomem_valid  (iomem_valid ),
		.iomem_ready  (iomem_ready ),
		.iomem_wstrb  (iomem_wstrb ),
		.iomem_addr   (iomem_addr  ),
		.iomem_wdata  (iomem_wdata ),
		.iomem_rdata  (iomem_rdata )
	);

/*
	assign debug_ser_tx = ser_tx;
	assign debug_ser_rx = ser_rx;

	assign debug_flash_csb = flash_csb;
	assign debug_flash_clk = flash_clk;
	assign debug_flash_io0 = flash_io0_di;
	assign debug_flash_io1 = flash_io1_di;
	assign debug_flash_io2 = flash_io2_di;
	assign debug_flash_io3 = flash_io3_di;
*/
endmodule
